`include "defines.svh"

import defines::*;

module app_mul_top(
	input sign,
	input scalar_t multiplicant,
	input scalar_t multiplier,
	output [63:0] product);
	
    logic [5:0] lod_multiplicant;
	logic [5:0] lod_multiplier;
	
	logic [30:0] frac_multiplicant;
	logic [30:0] frac_multiplier;
		
	logic [6:0] characteristic_sum;
	logic [31:0] fractional_sum_carry;
	logic [30:0] fractional_sum;
	logic [31:0] fractional_sum_corr_carry;
	logic [32:0] fractional_sum_appended;
	
	logic [94:0] internal_product;
	logic [46:0] shiftReg_multiplicant_tmp;
	logic [38:0] shiftReg_multiplicant;
    logic [46:0] shiftReg_multiplier_tmp;
    logic [38:0] shiftReg_multiplier;
	
	const logic [30:0] corr_factor = 30'b000101000000000000000000000000;
	
	assign product = internal_product[94:31];
	
	always_comb begin
            // Leading one detector for multiplicant 
            casez (multiplicant)
                32'b1???????????????????????????????: lod_multiplicant = 31;
                32'b01??????????????????????????????: lod_multiplicant = 30;
                32'b001?????????????????????????????: lod_multiplicant = 29;
                32'b0001????????????????????????????: lod_multiplicant = 28;
                32'b00001???????????????????????????: lod_multiplicant = 27;
                32'b000001??????????????????????????: lod_multiplicant = 26;
                32'b0000001?????????????????????????: lod_multiplicant = 25;
                32'b00000001????????????????????????: lod_multiplicant = 24;
                32'b000000001???????????????????????: lod_multiplicant = 23;
                32'b0000000001??????????????????????: lod_multiplicant = 22;
                32'b00000000001?????????????????????: lod_multiplicant = 21;
                32'b000000000001????????????????????: lod_multiplicant = 20;
                32'b0000000000001???????????????????: lod_multiplicant = 19;
                32'b00000000000001??????????????????: lod_multiplicant = 18;
                32'b000000000000001?????????????????: lod_multiplicant = 17;
                32'b0000000000000001????????????????: lod_multiplicant = 16;
                32'b00000000000000001???????????????: lod_multiplicant = 15;
                32'b000000000000000001??????????????: lod_multiplicant = 14;
                32'b0000000000000000001?????????????: lod_multiplicant = 13;
                32'b00000000000000000001????????????: lod_multiplicant = 12;
                32'b000000000000000000001???????????: lod_multiplicant = 11;
                32'b0000000000000000000001??????????: lod_multiplicant = 10;
                32'b00000000000000000000001?????????: lod_multiplicant = 9;
                32'b000000000000000000000001????????: lod_multiplicant = 8;
                32'b0000000000000000000000001???????: lod_multiplicant = 7;
                32'b00000000000000000000000001??????: lod_multiplicant = 6;
                32'b000000000000000000000000001?????: lod_multiplicant = 5;
                32'b0000000000000000000000000001????: lod_multiplicant = 4;
                32'b00000000000000000000000000001???: lod_multiplicant = 3;
                32'b000000000000000000000000000001??: lod_multiplicant = 2;
                32'b0000000000000000000000000000001?: lod_multiplicant = 1;
                32'b00000000000000000000000000000001: lod_multiplicant = 0;
                32'b00000000000000000000000000000000: lod_multiplicant = 0;
                default: lod_multiplicant = 0;
            endcase
                	
            // Leading one detector for multiplier.
            casez (multiplier)
                32'b1???????????????????????????????: lod_multiplier = 31;
                32'b01??????????????????????????????: lod_multiplier = 30;
                32'b001?????????????????????????????: lod_multiplier = 29;
                32'b0001????????????????????????????: lod_multiplier = 28;
                32'b00001???????????????????????????: lod_multiplier = 27;
                32'b000001??????????????????????????: lod_multiplier = 26;
                32'b0000001?????????????????????????: lod_multiplier = 25;
                32'b00000001????????????????????????: lod_multiplier = 24;
                32'b000000001???????????????????????: lod_multiplier = 23;
                32'b0000000001??????????????????????: lod_multiplier = 22;
                32'b00000000001?????????????????????: lod_multiplier = 21;
                32'b000000000001????????????????????: lod_multiplier = 20;
                32'b0000000000001???????????????????: lod_multiplier = 19;
                32'b00000000000001??????????????????: lod_multiplier = 18;
                32'b000000000000001?????????????????: lod_multiplier = 17;
                32'b0000000000000001????????????????: lod_multiplier = 16;
                32'b00000000000000001???????????????: lod_multiplier = 15;
                32'b000000000000000001??????????????: lod_multiplier = 14;
                32'b0000000000000000001?????????????: lod_multiplier = 13;
                32'b00000000000000000001????????????: lod_multiplier = 12;
                32'b000000000000000000001???????????: lod_multiplier = 11;
                32'b0000000000000000000001??????????: lod_multiplier = 10;
                32'b00000000000000000000001?????????: lod_multiplier = 9;
                32'b000000000000000000000001????????: lod_multiplier = 8;
                32'b0000000000000000000000001???????: lod_multiplier = 7;
                32'b00000000000000000000000001??????: lod_multiplier = 6;
                32'b000000000000000000000000001?????: lod_multiplier = 5;
                32'b0000000000000000000000000001????: lod_multiplier = 4;
                32'b00000000000000000000000000001???: lod_multiplier = 3;
                32'b000000000000000000000000000001??: lod_multiplier = 2;
                32'b0000000000000000000000000000001?: lod_multiplier = 1;
                32'b00000000000000000000000000000001: lod_multiplier = 0;
                32'b00000000000000000000000000000000: lod_multiplier = 0;
                default: lod_multiplier = 0;
            endcase



            // Barrel shifter for multiplicant's fractional part.
            shiftReg_multiplicant_tmp = {multiplicant, 31'b0} >> lod_multiplicant;
			shiftReg_multiplicant = shiftReg_multiplicant_tmp[38:0];
            frac_multiplicant = shiftReg_multiplicant[30:0];
		
	        // Barrel shifter for multipliers's fractional part.
		    shiftReg_multiplier_tmp = {multiplier, 31'b0} >> lod_multiplier;
		    shiftReg_multiplier = shiftReg_multiplier_tmp[38:0];
			frac_multiplier = shiftReg_multiplier[30:0];
	
            // Generate sum of fractional parts.
			fractional_sum_carry = {'0, frac_multiplicant} + {'0, frac_multiplier};
			fractional_sum = fractional_sum_carry[30:0];
			if(fractional_sum_carry[31]) begin
			     fractional_sum_corr_carry = {'0,fractional_sum} + ({'0,corr_factor} >> 1);
			     if (fractional_sum_corr_carry[31]) begin
			         fractional_sum_appended = { 2'b10, fractional_sum_corr_carry[30:0] };
			     end
			     else begin
                    fractional_sum_appended = { 2'b01, fractional_sum_corr_carry[30:0] };
			     end
			 end
			else begin
			     fractional_sum_corr_carry = {'0,fractional_sum} + {'0,corr_factor};
			     if (fractional_sum_corr_carry[31]) begin
			         fractional_sum_appended = { 2'b10, fractional_sum_corr_carry[30:0] };
			     end
			     else begin
                    fractional_sum_appended = { 2'b01, fractional_sum_corr_carry[30:0] };
			     end
			end
			
	        // Generate sum of characteristic parts.
			characteristic_sum = {'0,lod_multiplicant} + {'0,lod_multiplier} + {5'b0,fractional_sum_carry[31]};
	
            // Final barrel shifter.
            internal_product = {62'b0,fractional_sum_appended};
            internal_product = internal_product << characteristic_sum; 
            
            // Handle sign flag.
            // If signs of multiplier and multiplicant are unequal, the product has to be negative.
            // Therefore, the already calculated product, has to be negated (this equals to building
            // a 2-complement). 
            if(sign && (multiplicant[31] != multiplier[31])) begin
                internal_product = (~internal_product) + 1'b1; 
            end
        end
endmodule
